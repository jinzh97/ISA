module InstROM (
	input logic[9:0] InstAddress,
	output logic[8:0] InstOut
);

logic [8:0] rom [511:0];

assign InstOut = rom[InstAddress];

//Program 1
assign rom[0] = 'b000000000; //SETI 0
assign rom[1] = 'b110000000; //STORE 0 R0
assign rom[2] = 'b000011110; //SETI 30
assign rom[3] = 'b110000001; //STORE 0 R1
assign rom[4] = 'b101100000; //LOAD 0 R0
assign rom[5] = 'b011100001; //SEQ R1
assign rom[6] = 'b100010001; //BONE EXIT
assign rom[7] = 'b101110000; //LOAD 1 R0
assign rom[8] = 'b110001110; //STORE 0 R14
assign rom[9] = 'b101100000; //LOAD 0 R0
assign rom[10] = 'b001000001; //ADDI 1
assign rom[11] = 'b110000000; //STORE 0 R0
assign rom[12] = 'b101110000; //LOAD 1 R0
assign rom[13] = 'b110001111; //STORE 0 R15
assign rom[14] = 'b101101110; //LOAD 0 R14
assign rom[15] = 'b101000000; //PARITY 0
assign rom[16] = 'b110001100; //STORE 0 R12
assign rom[17] = 'b101101110; //LOAD 0 R14
assign rom[18] = 'b101000001; //PARITY 1
assign rom[19] = 'b110100001; //SHIFT 0 1
assign rom[20] = 'b010001100; //OR 0 R12
assign rom[21] = 'b110001100; //STORE 0 R12
assign rom[22] = 'b101101110; //LOAD 0 R14
assign rom[23] = 'b110100111; //SHIFT 0 7
assign rom[24] = 'b110110101; //SHIFT 1 5
assign rom[25] = 'b010001100; //OR 0 R12
assign rom[26] = 'b110001100; //STORE 0 R12
assign rom[27] = 'b101101110; //LOAD 0 R14
assign rom[28] = 'b101000010; //PARITY 2
assign rom[29] = 'b110100011; //SHIFT 0 3
assign rom[30] = 'b010001100; //OR 0 R12
assign rom[31] = 'b110001100; //STORE 0 R12
assign rom[32] = 'b101101110; //LOAD 0 R14
assign rom[33] = 'b110110001; //SHIFT 1 1
assign rom[34] = 'b110100101; //SHIFT 0 5
assign rom[35] = 'b110110001; //SHIFT 1 1
assign rom[36] = 'b010001100; //OR 0 R12
assign rom[37] = 'b110001100; //STORE 0 R12
assign rom[38] = 'b101101110; //LOAD 0 R14
assign rom[39] = 'b101000011; //PARITY 3
assign rom[40] = 'b110100111; //SHIFT 0 7
assign rom[41] = 'b010001100; //OR 0 R12
assign rom[42] = 'b110001100; //STORE 0 R12
assign rom[43] = 'b101101110; //LOAD 0 R14
assign rom[44] = 'b110110100; //SHIFT 1 4
assign rom[45] = 'b110001011; //STORE 0 R11
assign rom[46] = 'b101101111; //LOAD 0 R15
assign rom[47] = 'b110100100; //SHIFT 0 4
assign rom[48] = 'b010001011; //OR 0 R11
assign rom[49] = 'b110001011; //STORE 0 R11
assign rom[50] = 'b101100000; //LOAD 0 R0
assign rom[51] = 'b001011101; //ADDI 29
assign rom[52] = 'b110001010; //STORE 0 R10
assign rom[53] = 'b101101100; //LOAD 0 R12
assign rom[54] = 'b110011010; //STORE 1 R10
assign rom[55] = 'b101100000; //LOAD 0 R0
assign rom[56] = 'b001011110; //ADDI 30
assign rom[57] = 'b110001010; //STORE 0 R10
assign rom[58] = 'b101101011; //LOAD 0 R11
assign rom[59] = 'b110011010; //STORE 1 R10
assign rom[60] = 'b101100000; //LOAD 0 R0
assign rom[61] = 'b001000001; //ADDI 1
assign rom[62] = 'b110000000; //STORE 0 R0
assign rom[63] = 'b011010000; //JUMP LOOP
assign rom[64] = 'b111111111; //HALT


//program 2
assign rom[65] = 'b000010000; //SETI 10000
assign rom[66] = 'b110100010; //SHIFT 0 2
assign rom[67] = 'b110000000; //STORE 0 R0
assign rom[68] = 'b000011110; //SETI 11110
assign rom[69] = 'b010000000; //OR 0 R0
assign rom[70] = 'b110000001; //STORE 0 R1
assign rom[71] = 'b000001000; //SETI 8
assign rom[72] = 'b110000010; //STORE 0 R2
assign rom[73] = 'b101100000; //LOAD 0 R0 BEGINNING OF LOOP
assign rom[74] = 'b011100001; //SEQ R1
assign rom[75] = 'b100010010; //BONE EXIT
assign rom[76] = 'b101110000; //LOAD 1 R0
assign rom[77] = 'b110001110; //STORE 0 R14
assign rom[78] = 'b101100000; //LOAD 0 R0
assign rom[79] = 'b001000001; //ADDI 1
assign rom[80] = 'b110000000; //STORE 0 R0
assign rom[81] = 'b101110000; //LOAD 1 R0
assign rom[82] = 'b110001111; //STORE 0 R15
assign rom[83] = 'b101101110; //LOAD 0 R14
assign rom[84] = 'b110100110; //SHIFT 0 6
assign rom[85] = 'b110110110; //SHIFT 1 6
assign rom[86] = 'b110001100; //STORE 0 R12
assign rom[87] = 'b101101110; //LOAD 0 R14
assign rom[88] = 'b110100100; //SHIFT 0 4
assign rom[89] = 'b110110111; //SHIFT 1 7
assign rom[90] = 'b110100010; //SHIFT 0 2
assign rom[91] = 'b010001100; //OR 0 R12
assign rom[92] = 'b110001100; //STORE 0 R12
assign rom[93] = 'b101101110; //LOAD 0 R14
assign rom[94] = 'b110110111; //SHIFT 1 7
assign rom[95] = 'b110100011; //SHIFT 0 3
assign rom[96] = 'b010001100; //OR 0 R12
assign rom[97] = 'b110001100; //STORE 0 R12
assign rom[98] = 'b101101110; //LOAD 0 R14
assign rom[99] = 'b101000100; //PARITY 4
assign rom[100] = 'b110001011; //STORE 0 R11
assign rom[101] = 'b101101110; //LOAD 0 R14
assign rom[102] = 'b101000101; //PARITY 5
assign rom[103] = 'b110100001; //SHIFT 0 1
assign rom[104] = 'b010001011; //OR 0 R11
assign rom[105] = 'b110001011; //STORE 0 R11
assign rom[106] = 'b101101110; //LOAD 0 R14
assign rom[107] = 'b101000110; //PARITY 6
assign rom[108] = 'b110100010; //SHIFT 0 2
assign rom[109] = 'b010001011; //OR 0 R11
assign rom[110] = 'b110001011; //STORE 0 R11
assign rom[111] = 'b101101110; //LOAD 0 R14
assign rom[112] = 'b101000111; //PARITY 7
assign rom[113] = 'b110100011; //SHIFT 0 3
assign rom[114] = 'b010001011; //OR 0 R11
assign rom[115] = 'b110001011; //STORE 0 R11
assign rom[116] = 'b101101100; //LOAD 0 R12
assign rom[117] = 'b010011011; //OR 1 R11
assign rom[118] = 'b001100001; //SUBI 1
assign rom[119] = 'b110001010; //STORE 0 R10
assign rom[120] = 'b101100010; //LOAD 0 R2
assign rom[121] = 'b000101010; //SLT R10
assign rom[122] = 'b100010100; //BONE LOWER
assign rom[123] = 'b101101010; //LOAD 0 R10
assign rom[124] = 'b001101000; //SUBI 8
assign rom[125] = 'b110001010; //STORE 0 R10
assign rom[126] = 'b000000001; //SETI 1
assign rom[127] = 'b111001010; //SHIFTR 0 R10
assign rom[128] = 'b010011111; //OR 1 R15
assign rom[129] = 'b110001111; //STORE 0 R15
assign rom[130] = 'b011010101; //JUMP DECODE
assign rom[131] = 'b000000001; //SETI 1 BEGINNING OF LOWER
assign rom[132] = 'b111001010; //SHIFTR 0 R10
assign rom[133] = 'b010011110; //OR 1 R14
assign rom[134] = 'b110001110; //STORE 0 R14
assign rom[135] = 'b101101110; //LOAD 0 R14 BEGINNING OF DECODE
assign rom[136] = 'b110100101; //SHIFT 0 5 
assign rom[137] = 'b110110111; //SHIFT 1 7
assign rom[138] = 'b110001001; //STORE 0 R9
assign rom[139] = 'b101101110; //LOAD 0 R14
assign rom[140] = 'b110100001; //SHIFT 0 1 
assign rom[141] = 'b110110101; //SHIFT 1 5
assign rom[142] = 'b110100001; //SHIFT 0 1
assign rom[143] = 'b010001001; //OR 0 R9
assign rom[144] = 'b110001001; //STORE 0 R9
assign rom[145] = 'b101101111; //LOAD 0 R15
assign rom[146] = 'b110100100; //SHIFT 0 4
assign rom[147] = 'b010001001; //OR 0 R9
assign rom[148] = 'b110001001; //STORE 0 R9
assign rom[149] = 'b101101111; //LOAD 0 R15
assign rom[150] = 'b110110100; //SHIFT 1 4
assign rom[151] = 'b110001000; //STORE 0 R8
assign rom[152] = 'b101100000; //LOAD 0 R0
assign rom[153] = 'b001011101; //ADDI 29
assign rom[154] = 'b110001010; //STORE 0 R10
assign rom[155] = 'b101101001; //LOAD 0 R9
assign rom[156] = 'b110011010; //STORE 1 R10
assign rom[157] = 'b101100000; //LOAD 0 R0
assign rom[158] = 'b001011110; //ADDI 30
assign rom[159] = 'b110001010; //STORE 0 R10
assign rom[160] = 'b101101000; //LOAD 0 R8
assign rom[161] = 'b110011010; //STORE 1 R10
assign rom[162] = 'b101100000; //LOAD 0 R0
assign rom[163] = 'b001000001; //ADDI 1
assign rom[164] = 'b110000000; //STORE 0 R0
assign rom[165] = 'b011010011; //JUMP LOOP

//Program 3 PART 1
assign rom[166] = 'b000001010; //SETI 10
assign rom[167] = 'b110100100; //SHIFT 0 4
assign rom[168] = 'b110001101; //STORE 0 R13
assign rom[169] = 'b101111101; //LOAD 1 R13
assign rom[170] = 'b110001111; //STORE 0 R15
assign rom[171] = 'b000001000; //SETI 8
assign rom[172] = 'b110100100; //SHIFT 0 4
assign rom[173] = 'b110001110; //STORE 0 R14
assign rom[174] = 'b000000000; //SETI 0
assign rom[175] = 'b110000001; //STORE 0 R1
assign rom[176] = 'b110000000; //STORE 0 R0
assign rom[177] = 'b101101110; //LOAD 0 R14 //PART 1
assign rom[178] = 'b011101101; //SEQ R13
assign rom[179] = 'b100010110; //BONE PART2SETUP
assign rom[180] = 'b101111110; //LOAD 1 R14
assign rom[181] = 'b110110100; //SHIFT 1 4
assign rom[182] = 'b010011111; //OR 1 R15
assign rom[183] = 'b011100000; //SEQ R0
assign rom[184] = 'b010100001; //ADDR R1
assign rom[185] = 'b110000001; //STORE 0 R1
assign rom[186] = 'b101111110; //LOAD 1 R14
assign rom[187] = 'b110100001; //SHIFT 0 1
assign rom[188] = 'b110110100; //SHIFT 1 4
assign rom[189] = 'b010011111; //OR 1 R15
assign rom[190] = 'b011100000; //SEQ R0
assign rom[191] = 'b010100001; //ADDR R1
assign rom[192] = 'b110000001; //STORE 0 R1
assign rom[193] = 'b101111110; //LOAD 1 R14
assign rom[194] = 'b110100010; //SHIFT 0 2
assign rom[195] = 'b110110100; //SHIFT 1 4
assign rom[196] = 'b010011111; //OR 1 R15
assign rom[197] = 'b011100000; //SEQ R0
assign rom[198] = 'b010100001; //ADDR R1
assign rom[199] = 'b110000001; //STORE 0 R1
assign rom[200] = 'b101111110; //LOAD 1 R14
assign rom[201] = 'b110100011; //SHIFT 0 3
assign rom[202] = 'b110110100; //SHIFT 1 4
assign rom[203] = 'b010011111; //OR 1 R15
assign rom[204] = 'b011100000; //SEQ R0
assign rom[205] = 'b010100001; //ADDR R1
assign rom[206] = 'b110000001; //STORE 0 R1
assign rom[207] = 'b101111110; //LOAD 1 R14
assign rom[208] = 'b110100100; //SHIFT 0 4
assign rom[209] = 'b110110100; //SHIFT 1 4
assign rom[210] = 'b010011111; //OR 1 R15
assign rom[211] = 'b011100000; //SEQ R0
assign rom[212] = 'b010100001; //ADDR R1
assign rom[213] = 'b110000001; //STORE 0 R1
assign rom[214] = 'b101101110; //LOAD 0 R14
assign rom[215] = 'b001000001; //ADDI 1
assign rom[216] = 'b110001110; //STORE 0 R14
assign rom[217] = 'b011010111; //JUMP PART1
assign rom[218] = 'b000001100; //SETI 12 //PART2SETUP
assign rom[219] = 'b110100100; //SHIFT 0 4
assign rom[220] = 'b110000011; //STORE 0 R3
assign rom[221] = 'b101100001; //LOAD 0 R1
assign rom[222] = 'b110010011; //STORE 1 R3

//Program 3 PART 2
assign rom[223] = 'b000001000; //SETI 8
assign rom[224] = 'b110100100; //SHIFT 0 4
assign rom[225] = 'b110001110; //STORE 0 R14
assign rom[226] = 'b001000001; //ADDI 1
assign rom[227] = 'b110001100; //STORE 0 R12
assign rom[228] = 'b101101100; //LOAD 0 R12 //PART2
assign rom[229] = 'b011101101; //SEQ R13
assign rom[230] = 'b100011000; //BONE PART3SETUP
assign rom[231] = 'b101111110; //LOAD 1 R14
assign rom[232] = 'b110100101; //SHIFT 0 5
assign rom[233] = 'b110110100; //SHIFT 1 4
assign rom[234] = 'b110001011; //STORE 0 R11
assign rom[235] = 'b101111100; //LOAD 1 R12
assign rom[236] = 'b110110111; //SHIFT 1 7
assign rom[237] = 'b010001011; //OR 0 R11
assign rom[238] = 'b010011111; //OR 1 R15
assign rom[239] = 'b011100000; //SEQ R0
assign rom[240] = 'b010100001; //ADDR R1
assign rom[241] = 'b110000001; //STORE 0 R1
assign rom[242] = 'b101111110; //LOAD 1 R14
assign rom[243] = 'b110100110; //SHIFT 0 6
assign rom[244] = 'b110110100; //SHIFT 1 4
assign rom[245] = 'b110001011; //STORE 0 R11
assign rom[246] = 'b101111100; //LOAD 1 R12
assign rom[247] = 'b110110110; //SHIFT 1 6
assign rom[248] = 'b010001011; //OR 0 R11
assign rom[249] = 'b010011111; //OR 1 R15
assign rom[250] = 'b011100000; //SEQ R0
assign rom[251] = 'b010100001; //ADDR R1
assign rom[252] = 'b110000001; //STORE 0 R1
assign rom[253] = 'b101111110; //LOAD 1 R14
assign rom[254] = 'b110100111; //SHIFT 0 7
assign rom[255] = 'b110110100; //SHIFT 1 4
assign rom[256] = 'b110001011; //STORE 0 R11
assign rom[257] = 'b101111100; //LOAD 1 R12
assign rom[258] = 'b110110101; //SHIFT 1 5
assign rom[259] = 'b010001011; //OR 0 R11
assign rom[260] = 'b010011111; //OR 1 R15
assign rom[261] = 'b011100000; //SEQ R0
assign rom[262] = 'b010100001; //ADDR R1
assign rom[263] = 'b110000001; //STORE 0 R1
assign rom[264] = 'b101101110; //LOAD 0 R14
assign rom[265] = 'b001000001; //ADDI 1
assign rom[266] = 'b110001110; //STORE 0 R14
assign rom[267] = 'b001000001; //ADDI 1
assign rom[268] = 'b110001100; //STORE 0 R12
assign rom[269] = 'b011011001; //JUMP PART2
assign rom[270] = 'b101100011; //LOAD 0 R3 //PART3SETUP
assign rom[271] = 'b001000001; //ADDI 1
assign rom[272] = 'b110000011; //STORE 0 R3
assign rom[273] = 'b101100001; //LOAD 0 R1
assign rom[274] = 'b110010011; //STORE 1 R3

//Program 3 PART 3
assign rom[275] = 'b000000000; //SETI 0
assign rom[276] = 'b110000001; //STORE 0 R1
assign rom[277] = 'b000001000; //SETI 8
assign rom[278] = 'b110100100; //SHIFT 0 4
assign rom[279] = 'b110001110; //STORE 0 R14
assign rom[280] = 'b101101110; //LOAD 0 R14 //PART 3
assign rom[281] = 'b011101101; //SEQ R13
assign rom[282] = 'b100011010; //BONE EXIT
assign rom[283] = 'b101111110; //LOAD 1 R14
assign rom[284] = 'b110110100; //SHIFT 1 4
assign rom[285] = 'b010011111; //OR 1 R15
assign rom[286] = 'b011100000; //SEQ R0
assign rom[287] = 'b100011100; //BONE INC1
assign rom[288] = 'b101111110; //LOAD 1 R14
assign rom[289] = 'b110100001; //SHIFT 0 1
assign rom[290] = 'b110110100; //SHIFT 1 4
assign rom[291] = 'b010011111; //OR 1 R15
assign rom[292] = 'b011100000; //SEQ R0
assign rom[293] = 'b100011100; //BONE INC1
assign rom[294] = 'b101111110; //LOAD 1 R14
assign rom[295] = 'b110100010; //SHIFT 0 2
assign rom[296] = 'b110110100; //SHIFT 1 4
assign rom[297] = 'b010011111; //OR 1 R15
assign rom[298] = 'b011100000; //SEQ R0
assign rom[299] = 'b100011100; //BONE INC1
assign rom[300] = 'b101111110; //LOAD 1 R14
assign rom[301] = 'b110100011; //SHIFT 0 3
assign rom[302] = 'b110110100; //SHIFT 1 4
assign rom[303] = 'b010011111; //OR 1 R15
assign rom[304] = 'b011100000; //SEQ R0
assign rom[305] = 'b100011100; //BONE INC1
assign rom[306] = 'b101111110; //LOAD 1 R14
assign rom[307] = 'b110100100; //SHIFT 0 4
assign rom[308] = 'b110110100; //SHIFT 1 4
assign rom[309] = 'b010011111; //OR 1 R15
assign rom[310] = 'b011100000; //SEQ R0
assign rom[311] = 'b100111101; //BZERO INC2
assign rom[312] = 'b010100001; //ADDR R1 //INC
assign rom[313] = 'b110000001; //STORE 0 R1
assign rom[314] = 'b101101110; //LOAD 0 R14 //INC2
assign rom[315] = 'b001000001; //ADDI 1
assign rom[316] = 'b110001110; //STORE 0 R14
assign rom[317] = 'b011011011; //JUMP PART3
assign rom[318] = 'b101100011; //LOAD 0 R3 //EXIT
assign rom[319] = 'b001000001; //ADDI 1
assign rom[320] = 'b110000011; //STORE 0 R3
assign rom[321] = 'b101100001; //LOAD 0 R1
assign rom[322] = 'b110010011; //STORE 1 R3
assign rom[323] = 'b111111111; //EXIT

endmodule

